module my_or_gate (
    input wire A;
    input wire B;
    output wire OUT;
);

assign OUT = A | B // logical OR
    
endmodule